
module uart_testbench();
    reg clk_100mhz = 0; 
    reg clk_25mhz = 0;  
    reg rst=0;
    reg tx_start = 0;
    reg [7:0] tx_data = 8'hA5; 
    
    wire line;
    wire [7:0] rx_data;
    wire rx_done;
    wire tx_busy;

    
    always #5  clk_100mhz = ~clk_100mhz;
    always #20 clk_25mhz  = ~clk_25mhz; 
  reg [7:0]a;  
  
  
  
  transmitter transmitter_inst (
        .clk(clk_100mhz), 
        .reset(rst),          
        .data(tx_data),       
        .transmit(tx_start),  
        .txd(line),    
        .busy(tx_busy)  
    );

  
    receiver #(
        .clk_freq(25_000_000), 
      .baud_rate(9600)      
    ) receiver_inst (
        .clk_fpga(clk_25mhz), 
        .rst(rst),            
        .rxd(line),    
        .rxddata(rx_data),    
        .rdone(rx_done)      
    );
  
  initial begin 
    $dumpfile("testbench.vcd");
    $dumpvars(0,uart_testbench);
  end
  
    initial 
      begin
        $display("Starting");
        reset();
        send($random);
        check();
        #1000 
        $finish;
 end
  
  task reset; 
    begin 
   rst=1;
        #200 
      rst = 0;
    
  end 
  endtask
  task send( input [7:0]in);
    begin 
      wait(!tx_busy);
        @(posedge clk_100mhz);
        tx_start = 1;
        tx_data = in;
        a=in;
        @(posedge clk_100mhz);
        tx_start = 0;
  
  end
  endtask
  
  task check;
    begin
   fork
            begin
                wait(rx_done);
            end
            begin
                #2000000; 
                $display("Status: Timeout reached!");
            end
        join_any

    if (rx_data == a) begin
            $display("TEST PASSED");
        end else begin
          $display("TEST FAILED:  received %h , correct %h", rx_data,a);
        end
    end
  endtask
  
endmodule
